.title Ring Modulator
.include /home/gv/sys/fc14/fabrice/PySpice/examples/libraries/diode/standard-rectifier/1N4148.lib
Vmodulator in 0 DC 0V AC SIN(0V 1V 1000.0Hz 0s 0)
Vcarrier carrier 0 DC 0V AC SIN(0V 10V 100000.0Hz 0s 0)
Rin in 1 50
Linput 1 0 0.01
Linput_top input_top carrier 0.0025
Linput_bottom input_bottom carrier 0.0025
Kinput_top  Linput Linput_top 0.9
Kinput_bottom  Linput Linput_bottom 0.9
XD1 input_top output_top 1N4148
XD2 output_top input_bottom 1N4148
XD3 input_bottom output_bottom 1N4148
XD4 output_bottom input_top 1N4148
Loutput_top output_top 0 0.0025
Loutput_bottom output_bottom 0 0.0025
Loutput output 0 0.01
Koutput_top  Loutput Loutput_top 0.9
Koutput_bottom  Loutput Loutput_bottom 0.9
Rload output 0 1k
.options TNOM = 25
.options NOINIT
.options TEMP = 25
.options filetype = binary
* .ic V(output_bottom)=0 V(input_top)=0 V(input_bottom)=0 V(output_top)=0
.tran 5e-06 0.001
.end
