MOS OUTPUT CHARACTERISTICS
. OPTIONS NODE NOPAGE
VDS 3 0
VGS 2 0
M1 1 2 0 0 MOD1 L=4U W=6U AD=10P AS=10P
* VIDS MEASURES ID , WE COULD HAVE USED VDS, BUT ID WOULD BE NEGATIVE
VIDS 3 1
.MODEL MOD1 NMOS VTO=−2 NSUB= 1 . 0 E15 UO=550
. DC VDS 0 10 . 5 VGS 0 5 1
. END
